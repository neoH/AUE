// ******************************************************************************************
// File         : fetch_seqr.svh
// Author       : Ryan
// Creating Date: Thu Apr  2 20:13:48 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************
