// ******************************************************************************************
// File         : my_seqr.svh
// Author       : RyanHunter
// Creating Date: Sat May  2 06:59:07 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************


`ifndef my_seqr__svh
`define my_seqr__svh
`endif
