// ******************************************************************************************
// File         : fetcher_tb.sv
// Author       : RyanHunter
// Creating Date: Mon Apr  6 19:36:13 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************


`ifndef fetcher_tb__sv
`define fetcher_tb__sv

module fetcher_tb; // {





	initial begin // {
		run_test();
	end // }

endmodule // }

`endif
