// ******************************************************************************************
// File         : sce_dec_if.sv
// Author       : Ryan
// Creating Date: Tue Mar 31 22:15:52 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************

`ifndef sce_dec_if__sv
`define sce_dec_if__sv


interface sce_dec_if ;

	logic DEC2FET_VLD; // to fetch, valid



endinterface

`endif
