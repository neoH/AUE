// ******************************************************************************************
// File         : sce_define.sv
// Author       : Ryan
// Creating Date: Wed Apr  1 20:05:05 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************

`ifndef sce_define__sv
`define sce_define__sv



`endif
