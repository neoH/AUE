// ******************************************************************************************
// File         : my_dut.sv
// Author       : RyanHunter
// Creating Date: Sat May  2 06:58:59 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************


`ifndef my_dut__sv
`define my_dut__sv
`endif
