// ******************************************************************************************
// File         : head_import.svh
// Author       : Ryan
// Creating Date: Fri Apr  3 08:48:54 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************

`include "uvm_macros.svh"
import uvm_pkg::*;
import fetch_pkg::*;
