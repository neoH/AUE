// ******************************************************************************************
// File         : fetch_drv.svh
// Author       : Ryan
// Creating Date: Thu Apr  2 20:13:43 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************
