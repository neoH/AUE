// ******************************************************************************************
// File         : head_import.svh
// Author       : RyanHunter
// Creating Date: Tue Apr  7 09:06:23 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************


`ifndef head_import__svh
`define head_import__svh

`include "uvm_macros.svh"

import uvm_pkg::*;



`endif
