// ******************************************************************************************
// File         : fetch_rsp_item.svh
// Author       : Ryan
// Creating Date: Thu Apr  2 10:28:27 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************
