// ******************************************************************************************
// File         : rh_fu.sv
// Author       : RyanHunter
// Creating Date: Wed Apr 29 22:04:29 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************


`ifndef rh_fu__sv
`define rh_fu__sv


module RH_FU (
	fetch_mem_if.fetch fif,
	fetch_issue_if.fetch  iif
);





endmodule

`endif
