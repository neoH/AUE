// ******************************************************************************************
// File         : fetch_req_item.svh
// Author       : Ryan
// Creating Date: Thu Apr  2 10:28:21 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************

`ifndef fetch_req_item__svh
`define fetch_req_item__svh



`endif
