// ******************************************************************************************
// File         : tb_top.sv
// Author       : RyanHunter
// Creating Date: Wed Apr 22 09:57:13 2020
// Claim        : only the author can comment without a signature preffixed by ', that
// means anyone else want to change the code must comments with '.
// ******************************************************************************************


`ifndef tb_top__sv
`define tb_top__sv


`include "uvm_macros.svh"

module tb_top; // {

	import uvm_pkg::*;

	initial begin // {
		#1us;
		$finish;
	end // }


endmodule // }



`endif
